module CHECK1(
  input a, b,
  output f
);
  // Module Implementation

endmodule  // CHECK1