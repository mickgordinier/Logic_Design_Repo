// Declaring a new module with name 'Project05'
module Project05(
  input [16:0] SW,    // Using {SW[16], ..., SW[1], SW[0]} as inputs
  output [6:0] LEDR,  // Using {LEDR[6], ..., LEDR[0]} as outputs
  output [6:0] HEX0   // Using {HEX0[6], ..., HEX0[0]} as outputs
);
  // Module Implementation
  
endmodule  // Project 0.5