module Checker(
  input [6:0] A, B,
  output [6:0] F
);
  // Module Implementation

endmodule  // Checker